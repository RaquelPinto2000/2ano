---------------------------------------------------------------------------
-- University of Aveiro - DETI
-- "Computer Architecture I" course (Practical classes)
-- 
-- MIPS single-cycle datapath
---------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library work;
use work.DisplayUnit_pkg.all;
use work.MIPS_pkg.all;

entity MIPS_SingleCycle is
	port(	CLOCK_50 : in std_logic;
			KEY  		: in std_logic_vector(3 downto 0);
			SW   		: in std_logic_vector(17 downto 0);
			LEDR  	: out std_logic_vector(17 downto 0);
			LEDG  	: out std_logic_vector(8 downto 0);
			HEX0  	: out std_logic_vector(6 downto 0);
			HEX1  	: out std_logic_vector(6 downto 0);
			HEX2  	: out std_logic_vector(6 downto 0);
			HEX3  	: out std_logic_vector(6 downto 0);
			HEX4  	: out std_logic_vector(6 downto 0);
			HEX5  	: out std_logic_vector(6 downto 0);
			HEX6  	: out std_logic_vector(6 downto 0);
			HEX7  	: out std_logic_vector(6 downto 0));
end MIPS_SingleCycle;

architecture Shell of MIPS_SingleCycle is
-- Data signals
	signal sd_readData1 : std_logic_vector(31 downto 0);
	signal s_offset : std_logic_vector(31 downto 0);
-- Control signals (generated by the control unit)
	signal sc_RegDst : std_logic;

-- Signals related to the instruction code
	signal si_instr : std_logic_vector(31 downto 0);

-- Other signals
	signal s_clk : std_logic;
	signal s_pc : std_logic_vector(31 downto 0);
	
	signal s_rs : std_logic_vector(4 downto 0);
	signal s_rt : std_logic_vector(4 downto 0);
	signal s_rd : std_logic_vector(4 downto 0);
	signal s_mux1 : std_logic_vector(4 downto 0);
	signal s_mux2 : std_logic_vector(31 downto 0);
	signal s_alu : std_logic_vector(31 downto 0); -- sinal temporario
	signal s_readData1 : std_logic_vector(31 downto 0);
	signal s_readData2 : std_logic_vector(31 downto 0);
	signal s_funct : std_logic_vector(5 downto 0);
	signal s_AluControl:std_logic_vector(2 downto 0);
	signal s_opcode : std_logic_vector(5 downto 0);
	-- ControlUnit
	signal s_RegDst   :std_logic;
	signal s_Branch   :std_logic;
	signal s_Jump	   :std_logic;
	signal s_MemRead  :std_logic;
	signal s_MemWrite :std_logic;
	signal s_MemToReg :std_logic;
	signal s_ALUsrc   :std_logic;
	signal s_RegWrite :std_logic;
	signal s_ALUop : std_logic_vector(1 downto 0);
	--DataMemory
	signal s_readData : std_logic_vector(31 downto 0);
	signal s_mux3 : std_logic_vector(31 downto 0);
	
begin

-- PC Update
pcupd:	entity work.PCupdate(Behavioral)	
			port map(clk		=> s_clk,
						reset		=> not KEY(1),
						branch	=> '0',
						jump		=> '0',
						zero		=> '0',
						offset	=> s_offset,
						jAddr	=> sd_readData1(25 downto 0),
						pc			=> s_pc);

-- Instruction Memory
instmem:	entity work.InstructionMemory(Behavioral)
			generic map(ADDR_BUS_SIZE => ROM_ADDR_SIZE)
			port map(address		=> s_pc(7 downto 2),
						readData		=> sd_readData1);

-- Splitter
spliter:	entity work.InstrSplitter(Behavioral)
			port map(instruction		=> sd_readData1,
						opcode			=> s_opcode,
						rs					=> s_rs,
						rt					=> s_rt,
						rd					=> s_rd,
						funct				=> s_funct,
						imm				=> sd_readData1(15 downto 0),
						jAddr				=> sd_readData1(25 downto 0));
	
-- Sign Extender
signext:	entity work.SignExtend(Behavioral)
			port map(dataIn	=> sd_readData1(15 downto 0),
						dataOut	=> s_offset);
-- Mux1
mux1: entity work.Mux2N(Behavioral)
		generic map (N => 5)
		port map(sel => s_RegDst,
					input0 => s_rt,
					input1 => s_rd,
					muxout => s_mux1);
					
-- Mux2
mux2: entity work.Mux2N(Behavioral)
		generic map (N => 32)
		port map(sel => s_aLUsrc,
					input0 => s_readData2,
					input1 => s_offset,
					muxout => s_mux2);
--Mux3				
mux3: entity work.Mux2N(Behavioral)
		generic map (N => 32)
		port map(sel => s_memToReg,
					input0 => s_alu,
					input1 => s_readData,
					muxout => s_mux3);
					
-- Register file
regfile: entity work.RegFile(Strutural)
		port map (clk => s_clk,
					 writeEnable => sw(7),
					 writeReg  =>  s_mux1,
					 writeData  => s_mux3,  -- sinal temporario
					 readReg1 => s_rs,
					 readReg2  => s_rt,
					 readData1 => s_readData1,
					 readData2 => s_readData2);

-- Alucontrol
alucontrol: entity work.AluControlUnit( Behavioral)
	port map(ALUop => s_aLUop,
				funct => s_funct,
				ALUControl => s_AluControl);
-- ALU
alu: entity work.ALU32(Behavioral)
	port map (a => s_readData1,
				 b    => s_mux2,
				 oper => s_AluControl,
				 res  => s_alu, 
				 zero => open,
				 ovf => open);
				 
--	DU_RFdata <= s_instr;
--	DU_DMdata <= (s_alu);

dataMem: entity work.DataMemory(Behavioral)
	port map(clk       => s_clk, 
				readEn    => s_MemRead, 
				writeEn   => s_MemWrite, 
				address   => s_alu(7 downto 2), 
				writeData =>  s_readData2, 
				readData  => s_readData);
	
controlUnit: entity WORK.ControlUnit(Behavioral)
	port map( OpCode =>  s_opcode,
				RegDst =>  s_RegDst,
				Branch  =>  s_Branch,
				Jump	 =>s_Jump,
				MemRead => s_MemRead,
				MemWrite  => s_MemWrite,
				MemToReg  => s_MemToReg,
				ALUsrc    => s_ALUsrc,
				RegWrite  => s_RegWrite,
				ALUop     => s_ALUop);
				
LEDR(0)<=s_RegDst;
LEDR(1)<= s_Branch;
LEDR(2)<= s_Jump;
LEDR(3)<= s_MemRead;
LEDR(4) <= s_MemWrite;
LEDR(5) <= s_MemToReg;
LEDR(6) <= s_ALUsrc;
LEDR(7) <= s_RegWrite;
LEDR(9 downto 8) <= s_ALUop;
------------------------------------------------------------------------------
-- Support Modules						
------------------------------------------------------------------------------

-- Display Unit
display:	entity work.DisplayUnit(Behavioral)
			generic map(dataPathType => SINGLE_CYCLE_DP,
							IM_ADDR_SIZE => ROM_ADDR_SIZE,
							DM_ADDR_SIZE => RAM_ADDR_SIZE)
			port map(RefClk	=> CLOCK_50,
						InputSel	=> SW(1 downto 0),	
						DispMode	=> SW(17),
						NextAddr	=> KEY(3),
						Dir		=> KEY(2),
						disp0		=> HEX0,
						disp1		=> HEX1,
						disp2		=> HEX2,
						disp3		=> HEX3,
						disp4		=> HEX4,
						disp5		=> HEX5,
						disp6		=> HEX6,
						disp7		=> HEX7);		

-- Debouncer
debncer:	entity work.DebounceUnit(Behavioral)
			generic map(inPolarity	=> '0',
							outPolarity => '1')
			port map(refClk	=> CLOCK_50, 
						dirtyIn	=> KEY(0), 
						pulsedOut=> s_clk);						
end Shell;
